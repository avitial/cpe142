module dataMem();

endmodule
