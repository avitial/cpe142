module ctrlUnit();

endmodule
