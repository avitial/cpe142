module mux3to1();

endmodule
