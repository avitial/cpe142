module	fwdUnit();

endmodule
