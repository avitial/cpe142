module	hazDetnUnit();

endmodule
