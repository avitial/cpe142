/* Top Level */

'include “alu.v”
‘include “comptr.v”
‘include “ctrlUnit.v”  // still needs revision
‘include “dataMem.v”
‘include “fwdUnit.v”
‘include “hazDetnUnit.v”
‘include “instMem.v”
‘include “mux2to1.v”
‘include “opMux.v”
‘include “progCntr.v”
‘include “regDstDataMux.v”
‘include “regDstMux.v”
‘include “regFile.v”
‘include “signExtend.v”

module cpu(clk, rst);
	input clk, rst;

 




endmodule

