module fwdUnit();

endmodule
