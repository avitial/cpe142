module mux4to1();

endmodule
