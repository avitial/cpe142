module signExtend();

endmodule
