module dataMem(clk, rst, address, dataRead, dataWrite, MemRead, MemWrite);
  parameter addrSize = 16;
  parameter dataSize = 16;
  parameter Countloc = (1<< addrSize);

  input clk, rst;


endmodule
