module	dataMem();

endmodule
