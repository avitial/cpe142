module progrCntr();

endmodule
