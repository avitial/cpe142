module mux2to1();


endmodule
