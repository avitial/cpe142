'include "hazDetnUnit.v"
module

endmodule
