module comptr();

endmodule
