/* Top Level */

'include 

module 

endmodule
