module	instMem();

endmodule
