module mainCtrl();

endmodule
