'include "opMux.v"

module


endmodule
