module dataMem();
  parameter addrSize
  
endmodule
