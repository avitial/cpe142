module dataMem(clk, rst);
  parameter addrSize=16;
  parameter dataSize=16;
  


endmodule
